`timescale 1ns/1ns

module sonar_tb();